`ifndef _CFG_SVH_
`define _CFG_SVH_

`define RESETPC 32'h0000_0000

`endif /* !_CFG_SVH_ */
